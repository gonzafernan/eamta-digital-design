/*
 *  Module `signal_mux`
 *
 *  Generador y selector de se�ales.
 *
 *  Se generan las siguientes 4 se�ales con sus correspondientes archivos .hex:
 *  - Se�al 1: f1=1,5kHz y f2=17kHz (mem17khz.hex)
 *  - Se�al 2: f1=1,5kHz y f2=8,5kHz (mem17khz.hex)
 *  - Se�al 3: f1=1,5kHz y f2=5,66kHz (mem17khz.hex)
 *  - Se�al 4: f1=1,5kHz y f2=4,25kHz (mem17khz.hex)
 *  Luego dichas se�ales son entrada de un multiplexor que permite la seleccion
 *  de una de ellas segun i_sel[1:0].
 *
 *  Dependencias: modulo `signal_generator`
 *
 *  EAMTA 2021 - Digital Design
 *  Laboratorio 3: Integracion filtro FIR con memoria BRAM.
 *  Gonzalo G. Fernandez     10/03/2021
 *  File: signal_mux.v
 */

module signal_mux(
        i_clock,
        i_reset,
        i_sel,
        o_signal
    );

// Parameters
parameter NB_DATA   = 8;
parameter NB_COUNT  = 10;
parameter NB_SEL    = 2;

// Signals files
parameter MEM_SIG1_FILE = "D:\\digital_design_course\\eamta-digital-design\\lab3-fir_bram\\signals\\mem17khz.hex";
parameter MEM_SIG2_FILE = "D:\\digital_design_course\\eamta-digital-design\\lab3-fir_bram\\signals\\mem8p5khz.hex";
parameter MEM_SIG3_FILE = "D:\\digital_design_course\\eamta-digital-design\\lab3-fir_bram\\signals\\mem5p666khz.hex";
parameter MEM_SIG4_FILE = "D:\\digital_design_course\\eamta-digital-design\\lab3-fir_bram\\signals\\mem4p25khz.hex";

// Ports
input                               i_clock;
input                               i_reset;
input           [NB_SEL-1 : 0]      i_sel;
output  signed  [NB_DATA-1 : 0]     o_signal;

// Vars
reg     signed  [NB_DATA-1 : 0]     w_signal;   // mux output signal
wire    signed  [NB_DATA-1 : 0]     w_signal_1;
wire    signed  [NB_DATA-1 : 0]     w_signal_2;
wire    signed  [NB_DATA-1 : 0]     w_signal_3;
wire    signed  [NB_DATA-1 : 0]     w_signal_4;

// Signal 1 generation
signal_generator #
    (
    .NB_DATA(NB_DATA),
    .NB_COUNT(NB_COUNT),
    .MEM_INIT_FILE(MEM_SIG1_FILE)
    )
u_signal_gen_1
    (
    .i_clock(i_clock),
    .i_reset(i_reset), 
    .o_signal(w_signal_1)
    );

// Signal 2 generation
signal_generator #
    (
    .NB_DATA(NB_DATA),
    .NB_COUNT(NB_COUNT),
    .MEM_INIT_FILE(MEM_SIG2_FILE)
    )
u_signal_gen_2
    (
    .i_clock(i_clock),
    .i_reset(i_reset), 
    .o_signal(w_signal_2)
    );

// Signal 3 generation
signal_generator #
    (
    .NB_DATA(NB_DATA),
    .NB_COUNT(NB_COUNT),
    .MEM_INIT_FILE(MEM_SIG3_FILE)
    )
u_signal_gen_3
    (
    .i_clock(i_clock),
    .i_reset(i_reset), 
    .o_signal(w_signal_3)
    );

// Signal 4 generation
signal_generator #
    (
    .NB_DATA(NB_DATA),
    .NB_COUNT(NB_COUNT),
    .MEM_INIT_FILE(MEM_SIG4_FILE)
    )
u_signal_gen_4
    (
    .i_clock(i_clock),
    .i_reset(i_reset), 
    .o_signal(w_signal_4)
    );

// Multiplexer 4-to-1 (Language templates/Vivado)
always @(posedge i_clock) begin
    case (i_sel)
        2'b00: w_signal <= w_signal_1;
        2'b01: w_signal <= w_signal_2;
        2'b10: w_signal <= w_signal_3;
        2'b11: w_signal <= w_signal_4;
    endcase
end

assign o_signal = w_signal;

endmodule
